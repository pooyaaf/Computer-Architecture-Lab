module StageId(
 input clk, rst,
 input [31:0] PC,
 output [31:0] pcOut
);
endmodule